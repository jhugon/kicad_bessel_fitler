.title 7th Order LC circuit
r1 1 2 50
r2 100 0 50
c1 2 0 {C1:g}
l1 2 3 {L1:g}
c2 3 0 {C2:g}
l2 3 4 {L2:g}
c3 4 0 {C3:g}
l3 4 100 {L3:g}
c4 100 0 {C4:g}
.end
